library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity FullAdderNBits is
    generic (
        N : integer := 32  -- Número de bits
    );
    port (
        cin: in std_logic;
        x: in std_logic_vector(N-1 downto 0); 
        y: in std_logic_vector(N-1 downto 0);
        sigma: out std_logic_vector(N-1 downto 0);
        cout: out std_logic
    );
end entity FullAdderNBits;

architecture Structural of FullAdderNBits is
    component FullAdder
        port (
            cin: in std_logic;
            x: in std_logic;
            y: in std_logic;
            sigma: out std_logic;
            cout: out std_logic
        );
    end component;
    
    signal c: std_logic_vector(N downto 0); -- Acarreo interno
    
begin
    c(0) <= cin;
    
    generador: for i in 0 to N-1 generate
        FA: FullAdder port map (
            cin => c(i),
            x => x(i),
            y => y(i),
            sigma => sigma(i),
            cout => c(i+1)
        );
    end generate generador;
    
    cout <= c(N);

end Structural;
