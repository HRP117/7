library ieee;
use ieee.std_logic_1164.all;

entity FullAdder is
    port (
        cin: in std_logic;
        x: in std_logic;
        y: in std_logic;
        sigma: out std_logic;
        cout: out std_logic
    );
end entity FullAdder;

architecture DataFlow of FullAdder is
begin
    sigma <= cin xor x xor y;
    cout <= (cin and x) or (cin and y) or (x and y);
end DataFlow;
